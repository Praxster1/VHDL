library ieee;
use ieee.std_logic_1164.all;

package prng_pack is
    function min(a, b : integer) return integer;
    type polynom_array is array(natural range <>, natural range <>) of std_ulogic;

    constant prng_default_width : integer := 6;
    constant polynom_c : polynom_array(168 downto 1, 168 downto 1) :=
    (3 => (3 => '1', 2 => '1', others => '0'),
    4 => (4 => '1', 3 => '1', others => '0'),
    5 => (5 => '1', 3 => '1', others => '0'),
    6 => (6 => '1', 5 => '1', others => '0'),
    7 => (7 => '1', 6 => '1', others => '0'),
    8 => (8 => '1', 6 => '1', 5 => '1', 4 => '1', others => '0'),
    9 => (9 => '1', 5 => '1', others => '0'),
    10 => (10 => '1', 7 => '1', others => '0'),
    11 => (11 => '1', 9 => '1', others => '0'),
    12 => (12 => '1', 6 => '1', 4 => '1', 1 => '1', others => '0'),
    13 => (13 => '1', 4 => '1', 3 => '1', 1 => '1', others => '0'),
    14 => (14 => '1', 5 => '1', 3 => '1', 1 => '1', others => '0'),
    15 => (15 => '1', 14 => '1', others => '0'),
    16 => (16 => '1', 15 => '1', 13 => '1', 4 => '1', others => '0'),
    17 => (17 => '1', 14 => '1', others => '0'),
    18 => (18 => '1', 11 => '1', others => '0'),
    19 => (19 => '1', 6 => '1', 2 => '1', 1 => '1', others => '0'),
    20 => (20 => '1', 17 => '1', others => '0'),
    21 => (21 => '1', 19 => '1', others => '0'),
    22 => (22 => '1', 21 => '1', others => '0'),
    23 => (23 => '1', 18 => '1', others => '0'),
    24 => (24 => '1', 23 => '1', 22 => '1', 17 => '1', others => '0'),
    25 => (25 => '1', 22 => '1', others => '0'),
    26 => (26 => '1', 6 => '1', 2 => '1', 1 => '1', others => '0'),
    27 => (27 => '1', 5 => '1', 2 => '1', 1 => '1', others => '0'),
    28 => (28 => '1', 25 => '1', others => '0'),
    29 => (29 => '1', 27 => '1', others => '0'),
    30 => (30 => '1', 6 => '1', 4 => '1', 1 => '1', others => '0'),
    31 => (31 => '1', 28 => '1', others => '0'),
    32 => (32 => '1', 22 => '1', 2 => '1', 1 => '1', others => '0'),
    33 => (33 => '1', 2 => '1', others => '0'),
    34 => (34 => '1', 27 => '1', 2 => '1', 1 => '1', others => '0'),
    35 => (35 => '1', 33 => '1', others => '0'),
    36 => (36 => '1', 25 => '1', others => '0'),
    37 => (37 => '1', 5 => '1', 4 => '1', 3 => '1', 2 => '1', 1 => '1', others => '0'),
    38 => (38 => '1', 6 => '1', 5 => '1', 1 => '1', others => '0'),
    39 => (39 => '1', 35 => '1', others => '0'),
    40 => (40 => '1', 38 => '1', 21 => '1', 19 => '1', others => '0'),
    41 => (41 => '1', 38 => '1', others => '0'),
    42 => (42 => '1', 41 => '1', 20 => '1', 19 => '1', others => '0'),
    43 => (43 => '1', 42 => '1', 38 => '1', 37 => '1', others => '0'),
    44 => (44 => '1', 43 => '1', 18 => '1', 17 => '1', others => '0'),
    45 => (45 => '1', 44 => '1', 42 => '1', 41 => '1', others => '0'),
    46 => (46 => '1', 45 => '1', 26 => '1', 25 => '1', others => '0'),
    47 => (47 => '1', 42 => '1', others => '0'),
    48 => (48 => '1', 47 => '1', 21 => '1', 20 => '1', others => '0'),
    49 => (49 => '1', 4 => '1', others => '0'),
    50 => (50 => '1', 49 => '1', 24 => '1', 23 => '1', others => '0'),
    51 => (51 => '1', 50 => '1', 36 => '1', 35 => '1', others => '0'),
    52 => (52 => '1', 49 => '1', others => '0'),
    53 => (53 => '1', 52 => '1', 38 => '1', 37 => '1', others => '0'),
    54 => (54 => '1', 53 => '1', 18 => '1', 17 => '1', others => '0'),
    55 => (55 => '1', 31 => '1', others => '0'),
    56 => (56 => '1', 55 => '1', 35 => '1', 34 => '1', others => '0'),
    57 => (57 => '1', 5 => '1', others => '0'),
    58 => (58 => '1', 39 => '1', others => '0'),
    59 => (59 => '1', 58 => '1', 38 => '1', 37 => '1', others => '0'),
    60 => (60 => '1', 59 => '1', others => '0'),
    61 => (61 => '1', 60 => '1', 46 => '1', 45 => '1', others => '0'),
    62 => (62 => '1', 61 => '1', 6 => '1', 5 => '1', others => '0'),
    63 => (63 => '1', 62 => '1', others => '0'),
    64 => (64 => '1', 63 => '1', 61 => '1', 60 => '1', others => '0'),
    65 => (65 => '1', 47 => '1', others => '0'),
    66 => (66 => '1', 65 => '1', 57 => '1', 56 => '1', others => '0'),
    67 => (67 => '1', 66 => '1', 58 => '1', 57 => '1', others => '0'),
    68 => (68 => '1', 59 => '1', others => '0'),
    69 => (69 => '1', 67 => '1', 42 => '1', 40 => '1', others => '0'),
    70 => (70 => '1', 69 => '1', 55 => '1', 54 => '1', others => '0'),
    71 => (71 => '1', 65 => '1', others => '0'),
    72 => (72 => '1', 66 => '1', 25 => '1', 19 => '1', others => '0'),
    73 => (73 => '1', 48 => '1', others => '0'),
    74 => (74 => '1', 73 => '1', 59 => '1', 58 => '1', others => '0'),
    75 => (75 => '1', 74 => '1', 65 => '1', 64 => '1', others => '0'),
    76 => (76 => '1', 75 => '1', 41 => '1', 40 => '1', others => '0'),
    77 => (77 => '1', 76 => '1', 47 => '1', 46 => '1', others => '0'),
    78 => (78 => '1', 77 => '1', 59 => '1', 58 => '1', others => '0'),
    79 => (79 => '1', 7 => '1', others => '0'),
    80 => (80 => '1', 79 => '1', 43 => '1', 42 => '1', others => '0'),
    81 => (81 => '1', 77 => '1', others => '0'),
    82 => (82 => '1', 79 => '1', 47 => '1', 44 => '1', others => '0'),
    83 => (83 => '1', 82 => '1', 38 => '1', 37 => '1', others => '0'),
    84 => (84 => '1', 71 => '1', others => '0'),
    85 => (85 => '1', 84 => '1', 58 => '1', 57 => '1', others => '0'),
    86 => (86 => '1', 85 => '1', 74 => '1', 73 => '1', others => '0'),
    87 => (87 => '1', 74 => '1', others => '0'),
    88 => (88 => '1', 87 => '1', 17 => '1', 16 => '1', others => '0'),
    89 => (89 => '1', 51 => '1', others => '0'),
    90 => (90 => '1', 89 => '1', 72 => '1', 71 => '1', others => '0'),
    91 => (91 => '1', 90 => '1', 8 => '1', 7 => '1', others => '0'),
    92 => (92 => '1', 91 => '1', 80 => '1', 79 => '1', others => '0'),
    93 => (93 => '1', 91 => '1', others => '0'),
    94 => (94 => '1', 73 => '1', others => '0'),
    95 => (95 => '1', 84 => '1', others => '0'),
    96 => (96 => '1', 94 => '1', 49 => '1', 47 => '1', others => '0'),
    97 => (97 => '1', 91 => '1', others => '0'),
    98 => (98 => '1', 87 => '1', others => '0'),
    99 => (99 => '1', 97 => '1', 54 => '1', 52 => '1', others => '0'),
    100 => (100 => '1', 63 => '1', others => '0'),
    101 => (101 => '1', 100 => '1', 95 => '1', 94 => '1', others => '0'),
    102 => (102 => '1', 101 => '1', 36 => '1', 35 => '1', others => '0'),
    103 => (103 => '1', 94 => '1', others => '0'),
    104 => (104 => '1', 103 => '1', 94 => '1', 93 => '1', others => '0'),
    105 => (105 => '1', 89 => '1', others => '0'),
    106 => (106 => '1', 91 => '1', others => '0'),
    107 => (107 => '1', 105 => '1', 44 => '1', 42 => '1', others => '0'),
    108 => (108 => '1', 77 => '1', others => '0'),
    109 => (109 => '1', 108 => '1', 103 => '1', 102 => '1', others => '0'),
    110 => (110 => '1', 109 => '1', 98 => '1', 97 => '1', others => '0'),
    111 => (111 => '1', 101 => '1', others => '0'),
    112 => (112 => '1', 110 => '1', 69 => '1', 67 => '1', others => '0'),
    113 => (113 => '1', 101 => '1', others => '0'),
    114 => (114 => '1', 113 => '1', 57 => '1', 56 => '1', others => '0'),
    115 => (115 => '1', 114 => '1', 109 => '1', 107 => '1', others => '0'),
    116 => (116 => '1', 99 => '1', others => '0'),
    117 => (117 => '1', 116 => '1', 17 => '1', 16 => '1', others => '0'),
    118 => (118 => '1', 101 => '1', others => '0'),
    119 => (119 => '1', 118 => '1', 109 => '1', 108 => '1', others => '0'),
    120 => (120 => '1', 113 => '1', 9 => '1', 2 => '1', others => '0'),
    121 => (121 => '1', 103 => '1', others => '0'),
    122 => (122 => '1', 121 => '1', 63 => '1', 62 => '1', others => '0'),
    123 => (123 => '1', 121 => '1', others => '0'),
    124 => (124 => '1', 87 => '1', others => '0'),
    125 => (125 => '1', 124 => '1', 18 => '1', 17 => '1', others => '0'),
    126 => (126 => '1', 125 => '1', 90 => '1', 89 => '1', others => '0'),
    127 => (127 => '1', 126 => '1', others => '0'),
    128 => (128 => '1', 126 => '1', 101 => '1', 99 => '1', others => '0'),
    129 => (129 => '1', 124 => '1', others => '0'),
    130 => (130 => '1', 127 => '1', others => '0'),
    131 => (131 => '1', 130 => '1', 84 => '1', 83 => '1', others => '0'),
    132 => (132 => '1', 103 => '1', others => '0'),
    133 => (133 => '1', 132 => '1', 82 => '1', 81 => '1', others => '0'),
    134 => (134 => '1', 77 => '1', others => '0'),
    135 => (135 => '1', 124 => '1', others => '0'),
    136 => (136 => '1', 135 => '1', 11 => '1', 10 => '1', others => '0'),
    137 => (137 => '1', 116 => '1', others => '0'),
    138 => (138 => '1', 137 => '1', 131 => '1', 130 => '1', others => '0'),
    139 => (139 => '1', 136 => '1', 134 => '1', 131 => '1', others => '0'),
    140 => (140 => '1', 111 => '1', others => '0'),
    141 => (141 => '1', 140 => '1', 110 => '1', 109 => '1', others => '0'),
    142 => (142 => '1', 121 => '1', others => '0'),
    143 => (143 => '1', 142 => '1', 123 => '1', 122 => '1', others => '0'),
    144 => (144 => '1', 143 => '1', 75 => '1', 74 => '1', others => '0'),
    145 => (145 => '1', 93 => '1', others => '0'),
    146 => (146 => '1', 145 => '1', 87 => '1', 86 => '1', others => '0'),
    147 => (147 => '1', 146 => '1', 110 => '1', 109 => '1', others => '0'),
    148 => (148 => '1', 121 => '1', others => '0'),
    149 => (149 => '1', 148 => '1', 40 => '1', 39 => '1', others => '0'),
    150 => (150 => '1', 97 => '1', others => '0'),
    151 => (151 => '1', 148 => '1', others => '0'),
    152 => (152 => '1', 151 => '1', 87 => '1', 86 => '1', others => '0'),
    153 => (153 => '1', 152 => '1', others => '0'),
    154 => (154 => '1', 152 => '1', 27 => '1', 25 => '1', others => '0'),
    155 => (155 => '1', 154 => '1', 124 => '1', 123 => '1', others => '0'),
    156 => (156 => '1', 155 => '1', 41 => '1', 40 => '1', others => '0'),
    157 => (157 => '1', 156 => '1', 131 => '1', 130 => '1', others => '0'),
    158 => (158 => '1', 157 => '1', 132 => '1', 131 => '1', others => '0'),
    159 => (159 => '1', 128 => '1', others => '0'),
    160 => (160 => '1', 159 => '1', 142 => '1', 141 => '1', others => '0'),
    161 => (161 => '1', 143 => '1', others => '0'),
    162 => (162 => '1', 161 => '1', 75 => '1', 74 => '1', others => '0'),
    163 => (163 => '1', 162 => '1', 104 => '1', 103 => '1', others => '0'),
    164 => (164 => '1', 163 => '1', 151 => '1', 150 => '1', others => '0'),
    165 => (165 => '1', 164 => '1', 135 => '1', 134 => '1', others => '0'),
    166 => (166 => '1', 165 => '1', 128 => '1', 127 => '1', others => '0'),
    167 => (167 => '1', 161 => '1', others => '0'),
    168 => (168 => '1', 166 => '1', 153 => '1', 151 => '1', others => '0'),
    others => (others => '0')
    );

end prng_pack;

package body prng_pack is

    function min(a, b : integer) return integer is
    begin
        if a < b then
            return a;
        else
            return b;
        end if;
    end function min;

end package body;
