-------------------------------------------------------------------------------
-- Title      : sram controler - address path
-- Project    : 
-------------------------------------------------------------------------------
-- File       : sram_controler_address.vhd
-- Author     : Rabe
-- Company    : 
-- Created    : 2014-12-28
-- Last update: 2018-11-01
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2014 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-12-28  1.0      Rabe	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.sram_controler_pack.all;
entity sram_controler_address is

  port (
    clk_i : in std_ulogic;
    reset_n_i : in std_ulogic;
    fsm_we_i : in std_ulogic;
    fsm_re_i : in std_ulogic;
    fsm_start_addr_i : in std_ulogic_vector(18 downto 0);
    state_i : in FSM_T;
    srctr_end_addr_plus1_o : out std_ulogic_vector(18 downto 0);
    srctr_addr_reg_o : out std_ulogic_vector(18 downto 0));
end sram_controler_address;
architecture hehe of sram_controler_address is
  signal addr_reg : std_ulogic_vector(18 downto 0);
  signal addr_reg_plus1 : std_ulogic_vector(18 downto 0);
  --constant ONE : std_ulogic_vector(0 downto 0) := std_ulogic_vector(std_logic_vector(unsigned('1')());
begin


  addr_p : process (clk_i, reset_n_i)
  begin
    if reset_n_i = '1' then
      addr_reg <= (others => '1');
    elsif rising_edge(clk_i) then

      if (state_i = FSM_WRITE_MEM_33 or state_i = FSM_READ_MEM_33 or state_i = FSM_IDLE) and (fsm_re_i = '1' or fsm_we_i = '1') then
        srctr_addr_reg_o <= fsm_start_addr_i;
      elsif (state_i = FSM_WRITE_MEM_13 or state_i = FSM_WRITE_MEM_23 or state_i = FSM_READ_MEM_13 or state_i = FSM_READ_MEM_23) then
        addr_reg <= addr_reg_plus1;
      end if;
    end if;
  end process addr_p;

  adder_p : process (addr_reg)
  begin
    addr_reg_plus1 <= addr_reg + std_ulogic_vector(std_logic_vector(unsigned(1)));

  end process adder_p;

end architecture hehe;